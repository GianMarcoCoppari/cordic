LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;


PACKAGE CONFIG IS    
    CONSTANT M_BLOCKSIZE : INTEGER := 4; -- DIMENSIONE DI UN BLOCCO DI BIT
    CONSTANT M_BLOCKS    : INTEGER := 9; -- 36 BIT TOTALI
    CONSTANT M_BFRAC     : INTEGER := 7; -- 28 BIT FRAZIONARI
    
    CONSTANT PERIOD : TIME := 10 ns;
    CONSTANT M_CLA4LATENCY : INTEGER := 3; -- LATENZA DEL CLA4 IN COLPI DI CLOCK
    
    TYPE SUM_T IS RECORD 
        A   : STD_LOGIC_VECTOR(M_BLOCKSIZE * M_BLOCKS - 1 DOWNTO 0);
        B   : STD_LOGIC_VECTOR(M_BLOCKSIZE * M_BLOCKS - 1 DOWNTO 0);
        CIN : STD_LOGIC;
    END RECORD SUM_T;
    
    
END PACKAGE CONFIG;


PACKAGE BODY CONFIG IS 
END PACKAGE BODY CONFIG;
