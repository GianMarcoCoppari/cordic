LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
USE WORK.CONFIG.ALL;


PACKAGE CONFIGALU IS
    -- COSTANTI OPDOCE PER ALU.vhd
    -- Struttura OPCODE: 8 bit, 
    CONSTANT M_OPCODE_LENGTH : INTEGER := 8;
    
    -- MSB = 0: Op. Aritmetica, MSB = 1: Op. Logica
    CONSTANT M_LOGIC : STD_LOGIC := '0';
    CONSTANT M_ARITH : STD_LOGIC := '1';
    
    -- MSB - 1 = 0, Op. Unaria, MSB - 1 = 1, Op. Binaria
    CONSTANT M_UNARY  : STD_LOGIC := '0';
    CONSTANT M_BINARY : STD_LOGIC := '1';
    
    CONSTANT M_OPCODE_ADD  : STD_LOGIC_VECTOR(M_OPCODE_LENGTH - 1 DOWNTO 0) := M_ARITH & M_BINARY & "000000";
    CONSTANT M_OPCODE_SUB  : STD_LOGIC_VECTOR(M_OPCODE_LENGTH - 1 DOWNTO 0) := M_ARITH & M_BINARY & "000001";
    CONSTANT M_OPCODE_MULT : STD_LOGIC_VECTOR(M_OPCODE_LENGTH - 1 DOWNTO 0) := M_ARITH & M_BINARY & "000010";


END PACKAGE CONFIGALU;


PACKAGE BODY CONFIGALU IS 
END PACKAGE BODY CONFIGALU;