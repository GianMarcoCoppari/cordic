LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
USE WORK.CONFIG.ALL;


PACKAGE CONFIGCORDIC IS
    -- Constante per Numero di Iterazioni
    CONSTANT M_MAXITER : INTEGER := M_BLOCKSIZE * M_BFRAC;
    
    TYPE COORDS_T IS (M_CIRC, M_HYP);               -- Enumerazione per Tipo di Coordinate
    TYPE CORDICMODE_T IS (M_ROTATING, M_VECTORING); -- Enumerazione per Modalità di Lavoro
    
    
    TYPE LUT_T IS ARRAY (0 TO M_MAXITER - 1) OF STD_LOGIC_VECTOR(M_BLOCKSIZE * M_BLOCKS - 1 DOWNTO 0);
    CONSTANT M_ATANLUT : LUT_T := (
        X"000000000", X"000000000", X"000000000", X"000000000", 
        X"000000000", X"000000000", X"000000000", X"000000000", 
        X"000000000", X"000000000", X"000000000", X"000000000", 
        X"000000000", X"000000000", X"000000000", X"000000000", 
        X"000000000", X"000000000", X"000000000", X"000000000", 
        X"000000000", X"000000000", X"000000000", X"000000000", 
        X"000000000", X"000000000", X"000000000", X"000000000");
        
    CONSTANT NREP : INTEGER := 2;
    TYPE HINDEX_T IS ARRAY (0 TO M_MAXITER - 1 + NREP) OF INTEGER;
    CONSTANT M_HINDEX : HINDEX_T := (
        1, 2, 3, 4, 
        4, 5, 6, 7, 
        8, 9, 10, 11, 
        12, 13, 13, 14, 
        15, 16, 17, 18, 
        19, 20, 21, 22, 
        23, 24, 25, 26, 
        27, 28);
    
    CONSTANT M_ATANHLUT : LUT_T := (
        X"008C9F53D", X"004162BBE", X"00202B123", X"001005588", 
        X"000800AAC", X"000400155", X"00020002A", X"000100005", 
        X"000080000", X"000040000", X"000020000", X"000010000", 
        X"000008000", X"000004000", X"000002000", X"000001000", 
        X"000000800", X"000000400", X"000000200", X"000000100", 
        X"000000080", X"000000040", X"000000020", X"000000010", 
        X"000000008", X"000000004", X"000000002", X"000000001");
    
    
    -- Costanti di Configurazione per Algoritmo CORDIC
    TYPE CORDICSTATE_T IS RECORD 
        X : STD_LOGIC_VECTOR(M_BLOCKSIZE * M_BLOCKS - 1 DOWNTO 0);
        Y : STD_LOGIC_VECTOR(M_BLOCKSIZE * M_BLOCKS - 1 DOWNTO 0);
        Z : STD_LOGIC_VECTOR(M_BLOCKSIZE * M_BLOCKS - 1 DOWNTO 0);
    END RECORD;
    
    -- Costante (Inversa) di Guadagno
    CONSTANT M_KC : STD_LOGIC_VECTOR(M_BLOCKSIZE * M_BLOCKS - 1 DOWNTO 0) := X"000000000"; -- Circolare
    CONSTANT M_KY : STD_LOGIC_VECTOR(M_BLOCKSIZE * M_BLOCKS - 1 DOWNTO 0) := X"01351E872"; -- Iperbolico
   
    

    
    -- Costanti per la Riduzione del Range dell'Input
--    CONSTANT M_2PI : DATA_T := X"06487ED5";
--    CONSTANT M_PI2 : DATA_T := X"01921FB5";
--    CONSTANT M_LN2 : DATA_T := X"00B17217";
END PACKAGE CONFIGCORDIC;


PACKAGE BODY CONFIGCORDIC IS
END PACKAGE BODY CONFIGCORDIC;
